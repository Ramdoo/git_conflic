module moduleName (
    ports
);
    
    if () begin
        begin
        end
    end

    3333333
    3333333
    3333333
    2222222222222
    2222222222222
    2222222222222
    55555555555555
    55555555555555

endmodule