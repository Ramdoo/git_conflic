module moduleName (
    ports
);
    
    if () begin
        begin
        end
    end
endmodule