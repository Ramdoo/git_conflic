module moduleName (
    ports
);
    
    if () begin
        begin
        end
    end

    3333333
    3333333
    3333333
    2222222222222
    2222222222222
    2222222222222
    55555555555555
    55555555555555
    666666666666666
    777777777777
    888888888888
    888888888888
    999999999999
    1010

endmodule