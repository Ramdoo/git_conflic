module moduleName (
    ports
);
    
    if () begin
        begin
        end
    end

    2222222222222
    2222222222222
    2222222222222

endmodule