module moduleName (
    ports
);
    
    if () begin
        begin
        end
    end

    3333333
    3333333
    3333333

endmodule